../src/tt_um_theultimat_idli_top.v