`include "idli_pkg.svh"

// Top level of the core.
module idli_core_m import idli_pkg::*; (
  // Clock and reset.
  input  var logic          i_core_gck,
  input  var logic          i_core_rst_n,

  // SQI memory control interface.
  output var logic          o_core_sqi_sck,
  output var logic          o_core_sqi_cs,
  output var sqi_mode_t     o_core_sqi_mode,

  // SQI memory inputs and outputs.
  input  var logic  [3:0]   i_core_sqi_data,
  output var logic  [3:0]   o_core_sqi_data,

  // Data input interface.
  input  var logic  [3:0]   i_core_din,
  input  var logic          i_core_din_vld,
  output var logic          o_core_din_acp,

  // Data output interface.
  output var logic  [3:0]   o_core_dout,
  output var logic          o_core_dout_vld,
  input  var logic          i_core_dout_acp
);

  // {{{ Control Signals

  // Counter value and whether it's the final cycle.
  logic [1:0] ctr;
  logic       ctr_last_cycle;

  // }}} Control Signals

  // {{{ SQI Signals

  // Redirect signal as generated by the controller.
  logic sqi_redirect;

  // Data read from the SQI memory on this cycle.
  logic [3:0] sqi_rd_data;

  // }}} SQI Signals

  // {{{ Decode Signals

  // Whether data being presented to the decoder is valid.
  logic dcd_enc_vld;

  // Decoded instruction and whether it's valid.
  instr_t instr_q;
  instr_t instr_d;
  logic   instr_vld_q;

  // Whether the next instruction will take an immediate.
  logic dcd_next_instr_imm;

  // }}} Decode Signals

  // {{{ Register File Signals

  // General purpose register outputs.
  logic [3:0] grf_b_data;
  logic [3:0] grf_c_data;
  logic [3:0] grf_pc_data;

  // Predicate register outputs.
  logic prf_p_data;
  logic prf_q_data;

  // }}} Register File Signals

  // {{{ Execution Unit Signals

  // Whether the instruction should actually be executed.
  logic ex_instr_vld;

  // Outputs from the ALU.
  logic [3:0] alu_out;
  logic       alu_cout;

  // Operand C data input to the ALU and its source.
  logic [3:0] ex_op_c_data;
  logic       ex_op_c_imm;

  // }}} Execution Unit Signals


  // {{{ Control Logic

  idli_ctrl_m ctrl_u (
    .i_ctrl_gck             (i_core_gck),
    .i_ctrl_rst_n           (i_core_rst_n),

    .o_ctrl_ctr             (ctr),
    .o_ctrl_ctr_last_cycle  (ctr_last_cycle),

    .o_ctrl_sqi_redirect    (sqi_redirect),

    .i_ctrl_dcd_op_c_imm    (instr_d.op_c_imm),
    .o_ctrl_dcd_enc_vld     (dcd_enc_vld),

    .o_ctrl_ex_op_c_imm     (ex_op_c_imm)
  );

  // }}} Control Logic

  // {{{ SQI Logic

  idli_sqi_ctrl_m sqi_ctrl_u (
    .i_sqi_gck            (i_core_gck),
    .i_sqi_rst_n          (i_core_rst_n),

    .i_sqi_ctr            (ctr),
    .i_sqi_ctr_last_cycle (ctr_last_cycle),
    .i_sqi_redirect       (sqi_redirect),
    .i_sqi_rd             ('1),

    .o_sqi_sck            (o_core_sqi_sck),
    .o_sqi_cs             (o_core_sqi_cs),
    .o_sqi_mode           (o_core_sqi_mode),
    .i_sqi_rd_data        (i_core_sqi_data),
    .o_sqi_rd_data        (sqi_rd_data),
    .o_sqi_wr_data        (o_core_sqi_data),
    .i_sqi_wr_data        ('0),
    .i_sqi_wr_data_vld    ('1)
  );

  // }}} SQI Logic

  // {{{ Decode Logic

  idli_decode_m decode_u (
    .i_dcd_gck      (i_core_gck),
    .i_dcd_rst_n    (i_core_rst_n),

    .i_dcd_enc      (sqi_rd_data),
    .i_dcd_enc_vld  (dcd_enc_vld),

    .o_dcd_instr    (instr_d)
  );

  // Flop the decoded instruction once decoding is complete. Reset some of the
  // control signals that update state.
  always_ff @(posedge i_core_gck, negedge i_core_rst_n) begin
    if (!i_core_rst_n) begin
      instr_vld_q <= '0;
    end else if (ctr_last_cycle) begin
      instr_q     <= instr_d;
      instr_vld_q <= dcd_enc_vld;
    end
  end

  // Next instruction will take an immediate if the current instruction being
  // decoded indicates this, it's the last cycle, and the instruction in
  // decode is valid. We also make sure the current instruction executing is
  // valid as immediate data must come after a valid instruction has finished.
  always_comb dcd_next_instr_imm = dcd_enc_vld & ctr_last_cycle
                                 & instr_d.op_c_imm & instr_vld_q;

  // }}} Decode Logic

  // {{{ Register File Logic

  idli_grf_m grf_u (
    .i_grf_gck      (i_core_gck),

    .i_grf_b        (instr_q.op_b),
    .o_grf_b_data   (grf_b_data),

    .i_grf_c        (instr_q.op_c),
    .o_grf_c_data   (grf_c_data),

    .i_grf_a        (instr_q.op_a),
    .i_grf_a_vld    (instr_q.op_a_wr_en & ex_instr_vld),
    .i_grf_a_data   (alu_out),

    .i_grf_pc_vld   ('0),
    .i_grf_pc_data  ('x),
    .o_grf_pc_data  (grf_pc_data)
  );

  idli_prf_m prf_u (
    .i_prf_gck      (i_core_gck),

    .i_prf_p        (instr_q.op_p),
    .o_prf_p_data   (prf_p_data),

    .i_prf_q        (instr_q.op_q),
    .o_prf_q_data   (prf_q_data),
    .i_prf_q_wr_en  (instr_q.op_q_wr_en & ex_instr_vld),
    .i_prf_q_data   (alu_out[0])
  );

  // }}} Register File Logic

  // {{{ Execution Unit Logic

  idli_alu_m alu_u (
    .i_alu_gck    (i_core_gck),

    .i_alu_ctr_last_cycle (ctr_last_cycle),
    .i_alu_op             (instr_q.alu_op),

    .i_alu_lhs            (grf_b_data),
    .i_alu_rhs            (ex_op_c_data),

    .o_alu_out            (alu_out),
    .o_alu_cout           (alu_cout)
  );

  // Only actually execute an instruction if the predicate is non-zero.
  always_comb ex_instr_vld = prf_p_data & instr_vld_q;

  // Data for C comes from the GRF unless the control unit is indicating this
  // instruction takes immediate data - in this case the immediate used
  // directly from the memory.
  always_comb ex_op_c_data = ex_op_c_imm ? sqi_rd_data : grf_c_data;

  // }}} Execution Unit Logic

  // TODO Make use of the signals.
  logic _unused;

  always_comb o_core_din_acp     = '0;
  always_comb o_core_dout        = '0;
  always_comb o_core_dout_vld    = '0;

  always_comb _unused = &{i_core_din, i_core_dout_acp, i_core_din_vld, 1'b0,
    prf_p_data, prf_q_data, alu_cout};

endmodule
